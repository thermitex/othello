module othello(
    
);

endmodule // othello